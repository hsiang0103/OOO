`include "riscv_instr_gen_config_ext.sv"