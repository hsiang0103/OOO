// program start address
`define RESET_ADDR 32'h0000_2000

// Issue Queue
`define IQ_LEN      16

// Load Queue
`define LQ_LEN      16

// Store Queue
`define SQ_LEN      16

// Reorder Buffer
`define ROB_LEN     16

// Inst Queue
`define INST_QUEUE_LEN 4