// program start address
`define RESET_ADDR 32'h0000_2000

// Issue Queue
`define IQ_LEN      4

// Load Queue
`define LQ_LEN      4

// Store Queue
`define SQ_LEN      4

// Reorder Buffer
`define ROB_LEN     8